module top_module(
    output zero
);
    assign zero = 0;// Module body starts after semicolon

endmodule
